module decoder198 (a, b, c, d, e, f, g, h, a0, b0, c0, d0, e0, f0, g0, a10, b10, c10, d10, e10, f10, g10, a20, b20, c20, d20, e20, f20, g20);
	input a, b, c, d, e, f, g, h;
	output a0, b0, c0, d0, e0, f0, g0, a10, b10, c10, d10, e10, f10, g10, a20, b20, c20, d20, e20, f20, g20;
	assign a0 = ((a) | (b&c&f) | | (b&c&e) | (b&c&d));
	assign b0 = 0;
	assign c0 = 0;
	assign d0 = ((a) | (b&c&f) | | (b&c&e) | (b&c&d));
	assign e0 = ((a) | (b&c&f) | | (b&c&e) | (b&c&d));
	assign f0 = ((a) | (b&c&f) | | (b&c&e) | (b&c&d));
	assign g0 = 1;
	
	assign a10 = ((b&c&d&~e) | (~a&~b&~d&e&g) | (~b&~c&~d&e&f) | (~b&~c&d&~e&~f) | (~a&~b&c&~d&e) | (a&~c&d&~e&~g) | (~a&~b&d&~e&~f&~g) | (~a&c&~d&e&f&g));
	assign b10 = ((a&~c&d&e) | (a&c&~d&~e) | (~a&~b&c&d&g) | (~a&~b&c&d&f) | (~a&~b&c&d&e) | (a&~c&d&f&g) | (a&c&~d&~f&~g) | (~a&b&~c&~d&~e&~f) | (~a&b&~c&~d&~e&~g));
	assign c10 = ((b&c&d&e) | (~a&~b&~c&d&~e&f) | (~a&~b&~c&d&f&~g) | (~a&~b&~c&d&e&~f) | (a&~b&~c&~d&~e&~f&~g));
	assign d10 = ((~b&~d&e&f) | (~d&e&f&g) | (b&~c&~d&e) | (b&c&d&~e) | (a&d&~e&~f) | (~a&~b&~d&e&g) | (~b&~c&d&~e&~f) | (~b&d&~e&~f&~g) | (~a&~b&c&~d&e) | (~b&c&~d&e&g) | (a&~c&d&~e&~g) | (~a&b&~c&~d&f&g));
	assign e10 = ((a&b) | (a&~c&g) | (a&~c&f) | (a&~c&e) | (~b&~d&e&g) | (~b&~d&e&f) | (~b&d&~e&~f) | (~a&~b&c&~d) | (~a&~b&c&~f) | (~a&c&~e&~f) | (~a&c&d&~e) | (~c&e&f&g) | (~d&e&f&g) | (b&~c&~d&e) | (b&~c&e&g) | (b&~c&e&f) | (a&e&f&g) | (b&~c&~d&f&g));
	assign f10 = ((b&c&d) | (~a&~b&~c&d) | (b&~c&~d&e) | (~a&~b&~c&e&g) | (~a&~b&~c&e&f) | (~a&~b&c&~d&~e) | (a&~b&~c&~d&~e) | (a&~b&~c&~d&~f) | (b&~d&e&f&g) | (a&~d&e&~f&g) | (a&c&~d&e&f) | (a&c&d&~e&~f) | (~a&b&~c&~d&f&g));
	assign g10 = ((b&~d&e) | (~a&~b&~c&~d) | (b&c&~d&f) | (b&c&d&~e) | (~a&~b&~c&~e&~f) | (~a&~c&~d&f&g) | (a&c&~d&e&g) | (a&c&~d&e&f) | (a&c&d&~e&~f));
	
	assign a20 = ((a&b&~f&g&~h) | (b&~c&~d&~e&f&g&h) | (b&~c&~d&e&~f&g&~h) | (b&~c&d&~e&~f&~g&h) | (b&~c&d&~e&f&~g&~h) | (b&~c&d&e&~f&g&h) | (b&~c&d&e&f&g&~h) | (b&c&~d&~e&f&~g&h) | (b&c&~d&e&~f&~g&~h) | (b&c&~d&e&f&g&h) | (b&c&d&~e&~f&g&~h) | (b&c&d&e&~f&~g&h) | (b&c&d&e&f&~g&~h) | (a&~c&~d&e&f&~g&h) | (a&~c&d&~e&~f&~g&~h) | (a&~c&d&~e&f&g&h) | (a&~c&d&e&~f&g&~h) | (a&c&~d&~e&~f&~g&h) | (a&c&~d&~e&f&~g&~h) | (a&c&~d&e&~f&g&h) | (a&c&~d&e&f&g&~h) | (a&c&d&~e&f&~g&h) | (a&c&d&e&~f&~g&~h) | (a&c&d&e&f&g&h) | (~a&~b&~c&~d&~e&~f&~g&h) | (~a&~b&~c&~d&~e&f&~g&~h) | (~a&~b&~c&~d&e&~f&g&h) | (~a&~b&~c&~d&e&f&g&~h) | (~a&~b&~c&d&~e&f&~g&h) | (~a&~b&~c&d&e&~f&~g&~h) | (~a&~b&~c&d&e&f&g&h) | (~a&~b&c&~d&~e&~f&g&~h) | (~a&~b&c&~d&e&~f&~g&h) | (~a&~b&c&~d&e&f&~g&~h) | (~a&~b&c&d&~e&~f&g&h) | (~a&~b&c&d&~e&f&g&~h) | (~a&~b&c&d&e&f&~g&h) | (~a&b&~c&~d&~e&~f&~g&~h) | (a&~b&~c&~d&~e&~f&g&h) | (a&~b&~c&~d&~e&f&g&~h));
	assign b20 = ((a&b&g&h) | (a&b&f&~g&~h) | (b&~c&~d&e&~f&g&h) | (b&~c&~d&e&f&~g&~h) | (b&~c&d&~e&f&~g&h) | (b&~c&d&~e&f&g&~h) | (b&~c&d&e&f&g&h) | (b&c&~d&~e&~f&~g&~h) | (b&c&~d&e&~f&~g&h) | (b&c&~d&e&~f&g&~h) | (b&c&d&~e&~f&g&h) | (b&c&d&~e&f&~g&~h) | (b&c&d&e&f&~g&h) | (b&c&d&e&f&g&~h) | (a&~c&~d&~e&f&g&h) | (a&~c&~d&e&~f&~g&~h) | (a&~c&d&~e&~f&~g&h) | (a&~c&d&~e&~f&g&~h) | (a&~c&d&e&~f&g&h) | (a&~c&d&e&f&~g&~h) | (a&c&~d&~e&f&~g&h) | (a&c&~d&~e&f&g&~h) | (a&c&~d&e&f&g&h) | (a&~c&~d&e&~f&~g&~h) | (a&c&d&~e&~f&~g&~h) | (a&c&d&e&~f&~g&h) | (a&c&d&e&~f&g&~h) | (~a&~b&~c&~d&~e&f&~g&h) | (~a&~b&~c&~d&~e&f&g&~h) | (~a&~b&~c&~d&e&f&g&h) | (~a&~b&~c&d&~e&~f&~g&~h) | (~a&~b&~c&d&e&~f&~g&h) | (~a&~b&~c&d&e&~f&g&~h) | (~a&~b&c&~d&~e&~f&g&h) | (~a&~b&c&~d&~e&f&~g&~h) | (~a&~b&c&~d&e&f&~g&h) | (~a&~b&c&~d&e&f&g&~h) | (~a&~b&c&d&~e&f&g&h) | (~a&~b&c&d&e&~f&~g&~h) | (~a&b&~c&~d&~e&~f&~g&h) | (~a&b&~c&~d&~e&~f&g&~h));
	assign c20 = ((a&b&~f&~g&~h) | (b&~c&~d&e&~f&~g&~h) | (b&~c&d&~e&~f&g&~h) | (b&~c&d&e&f&~g&~h) | (b&c&~d&~e&f&g&~h) | (b&c&d&~e&~f&~g&~h) | (b&c&d&e&~f&g&~h) | (b&~c&~d&e&~f&~g&~h) | (a&~c&~d&e&f&g&~h) | (a&~c&d&e&~f&~g&~h) | (a&c&~d&~e&~f&g&~h) | (a&c&~d&e&f&~g&~h) | (a&c&d&~e&f&g&~h) | (~a&~b&~c&~d&~e&~f&g&~h) | (~a&~b&~c&~d&e&f&~g&~h) | (~a&~b&~c&d&~e&f&g&~h) | (~a&~b&c&~d&~e&~f&~g&~h) | (~a&~b&c&~d&e&~f&g&~h) | (~a&~b&c&d&~e&f&~g&~h) | (~a&~b&c&d&e&f&g&~h) | (a&~b&~c&~d&~e&f&~g&~h));
	assign d20 = ((a&b&f&h) | (a&b&~f&g&~h) | (b&~c&~e&f&g&h) | (b&c&~d&~e&~g&h) | (b&c&~e&f&~g&h) | (b&c&~d&e&g&h) | (b&c&e&f&g&h) | (a&~c&~d&e&~g&h) | (a&~c&e&f&~g&h) | (a&~c&d&~e&g&h) | (a&c&~e&~f&~g&h) | (a&c&e&~f&g&h) | (a&c&d&~e&~g&h) | (a&c&d&e&g&h) | (~a&~b&~c&~f&~e&~g&h) | (~a&~c&~d&~e&f&g&h)  | (~a&~b&~c&e&~f&g&h) | (~a&~b&~c&d&~e&~g&h) | (~a&~c&d&~e&~f&~g&h) | (~a&~b&~c&d&e&g&h) | (~a&~c&d&e&~f&g&h) | (~a&c&~d&~e&f&~g&h) | (~a&~b&c&e&~f&~g&h) | (~a&c&~d&e&f&g&h) | (~a&~b&c&d&e&~g&h) | (~a&c&d&e&~f&~g&h) | (~a&b&~c&~d&~e&g&h) | (a&~b&~c&~e&~f&g&h) | (b&~c&~d&e&~f&g&~h) | (b&~c&~d&e&f&~g&h) | (b&~c&d&~e&f&~g&~h) | (b&~c&d&e&f&g&~h) | (b&c&~d&e&~f&~g&~h) | (b&c&d&~e&~f&g&~h) | (b&c&d&e&f&~g&~h) | (a&~c&d&~e&~f&~g&~h) | (a&~c&d&e&~f&g&~h) | (a&c&~d&~e&f&~g&~h) | (a&c&~d&~e&f&g&h) | (a&c&~d&e&f&g&~h) | (a&c&d&e&~f&~g&~h) | (~a&~b&~c&~d&~e&f&~g&~h) | (~a&~b&~c&~d&e&f&g&~h) | (~a&~b&~c&d&e&~f&~g&~h) | (~a&~b&c&~d&~e&~f&g&~h) | (~a&~b&c&~d&e&f&~g&~h) | (~a&~b&c&d&~e&~f&g&h) | (~a&~b&c&d&~e&f&g&~h) | (a&~b&~c&~d&~e&f&g&~h) | (~a&b&~c&~d&~e&~f&~g&~h));      
	assign e20 = ((h) | (a&b&~f&g) | (b&~c&~d&e&~f&g) | (b&~c&d&~e&f&~g) | (b&~c&d&e&f&g) | (b&c&~d&e&~f&~g) | (b&c&d&~e&~f&g) | (b&c&d&e&f&~g) | (a&~c&d&~e&~f&~g) | (a&~c&d&e&~f&g) | (a&c&~d&~e&f&~g) | (a&c&~d&e&f&g) | (a&c&d&e&~f&~g) | (~a&~b&~c&~d&~e&f&~g) | (~a&~b&~c&~d&e&f&g) | (~a&~b&~c&d&e&~f&~g) | (~a&~b&c&~d&~e&~f&g) | (~a&~b&c&~d&e&f&~g) | (~a&~b&c&d&~e&f&g) | (~a&b&~c&~d&~e&~f&~g) | (a&~b&~c&~d&~e&f&g));
	assign f20 = ((a&b&~f&~g) | (a&b&~g&h) | (a&~c&e&~g&h) | (~a&~c&~d&~e&g&h) | (~a&~c&~d&~e&g&h) | (~a&~c&~e&f&g&h) | (~a&c&~d&~e&~g&h) | (~a&c&~d&e&g&h) | (~c&~d&e&f&~g&h) | (c&d&~e&f&~g&h) | (c&d&e&f&g&h) | (b&~c&~d&e&~f&~g) | (b&~c&d&~e&~f&h) | (b&~c&d&~e&~f&g) | (b&~c&d&~f&g&h) | (b&~c&d&e&f&~g) | (b&c&~d&~e&f&g) | (b&c&d&~e&~f&~g) | (b&c&d&~f&~g&h) | (b&c&d&e&~f&g) | (a&~c&~d&e&f&g) | (a&~c&d&~e&g&h) | (a&~c&d&e&~f&~g) | (a&c&~e&~f&~g&h) | (a&c&~d&~e&~f&g) | (a&c&~d&~e&g&h) | (a&c&e&~f&g&h) | (a&c&~d&e&f&~g) | (a&c&d&~e&f&g) | (~a&~b&~c&~d&~e&~f&h) | (~a&~b&~c&~d&~e&~f&g) | (~b&~c&~d&~e&~f&g&h) | (~a&~b&~c&e&~f&g&h) | (~a&~b&~c&~d&e&f&~g) | (~a&~b&~c&d&~e&~g&h) | (~a&~b&~c&d&~e&f&g) | (~a&~b&~c&d&f&g&h) | (~a&~b&c&~d&~e&~f&~g) | (~a&~b&c&e&~f&~g&h) | (~a&~b&c&~d&e&~f&g) | (~a&~b&c&d&~e&f&~g) | (~a&~b&c&d&f&~g&h) | (~a&~b&c&d&e&f&g) | (a&~b&~c&~d&~e&f&~g) | (~a&~b&c&d&~e&~f&g&h));
	assign g20 = ((a&b&f&h) | (b&~c&~e&f&g&h) | (b&~c&d&~e&~f&~g) | (b&~c&d&e&~f&g) | (b&c&~d&~e&~g&h) | (b&c&~d&~e&f&~g) | (b&c&~e&f&~g&h) | (b&c&~d&e&g&h) | (b&c&~d&e&f&g) | (b&c&e&f&g&h) | (b&c&d&e&~f&~g) | (a&~c&~d&e&~g&h) | (a&~c&~d&e&f&~g) | (a&~c&e&f&~g&h) | (a&~c&d&~e&g&h) | (a&~c&d&~e&f&g) | (a&c&~d&~e&~f&~g) | (a&c&~e&~f&~g&h) | (a&c&~d&e&~f&g) | (a&c&e&~f&g&h) | (a&c&d&~e&f&~g) | (a&c&d&e&f&g) | (~a&~b&~c&~d&~e&~f&~g) | (~a&~b&~c&~e&~f&~g&h) | (~a&~c&~d&~e&f&g&h) | (~a&~b&~c&~d&e&~f&g) | (~a&~b&~c&e&~f&g&h) | (~a&~b&~c&d&~e&f&~g) | (~a&~b&~c&d&e&f&g) | (~a&c&~d&~e&f&~g&h) | (~a&~b&c&~d&e&~f&~g) | (~a&~b&c&e&~f&~g&h) | (~a&c&~d&e&f&g&h) | (~a&~b&c&d&~e&~f&g) | (~a&~b&c&d&e&f&~g) | (~a&b&~c&~d&~e&g&h) | (~a&b&~c&~d&~e&f&g) | (a&~b&~c&~d&~e&~f&g) | (b&~c&~d&e&f&~g&h) | (a&c&~d&~e&f&g&h));
endmodule
