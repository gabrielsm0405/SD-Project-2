module decoder99 (e0, e1, e2, e3, e4, e5, e6, a, b, c, d, e, f, g, a10, b10, c10, d10, e10, f10, g10);
	input e0, e1, e2, e3, e4, e5, e6;
	output a, b, c, d, e, f, g, a10, b10, c10, d10, e10, f10, g10;
	
	assign a = ((e1&~e2&e3) | (~e0&~e2&e3&e5) | (~e0&~e2&e3&e4) | (~e0&~e1&e2&~e3&~e4) | (~e0&e2&~e3&~e4&~e5));
	assign b = ((e1&e2&e5) | (e1&e2&e4) | (e1&e2&e3) | (e0&~e1&~e2&~e3&~e4) | (e0&~e1&~e2&~e3&~e5));
	assign c = ((~e0&~e1&e2&~e3&e4) | (~e0&~e1&e2&e4&~e5) | (~e0&~e1&e2&e3&~e4));
	assign d = ((~e2&e3&e5) | (~e2&e3&e4) | (~e2&e3&e1) | (~e2&e3&e0) | (e0&~e2&e4&e5) | (~e0&~e1&e2&~e3&~e4) | (~e0&~e5&e2&~e3&~e4));
	assign e = ((e1&~e3) | (e1&~e4) | (~e2&e3&e5) | (~e2&e3&e4) | (~e2&e0&e3) | (e0&e3&e5) | (e0&e3&e4) | (~e1&e3&e4&e5) | (~e0&e2&~e3&~e4) | (e0&~e2&e4&e5));
	assign f = ((~e0&~e1&e2) | (e0&~e2&e3) | (~e0&~e1&e3&e5) | (~e0&~e1&e3&e4) | (~e0&e1&~e2&~e3) | (e0&~e2&e4&e5));
	assign g = ((~e0&~e1&~e2) | (e3&~e1&~e2) | (~e0&~e1&~e3&~e4) | (~e1&~e2&e4&e5));  
	assign a10 = ((e1&~e2&e3&~e4&~e5&e6) | (e1&~e2&e3&e4&~e5&~e6) | (e1&e2&~e3&~e4&e5&e6) | (e1&e2&~e3&e4&e5&~e6) | (e1&e2&e3&e4&~e5&e6) | (e0&~e2&~e3&e4&e5&e6) | (e0&~e2&e3&~e4&e5&~e6) | (e0&e2&~e3&~e4&~e5&e6) | (e0&e2&~e3&e4&~e5&~e6) | (e0&e2&e3&~e4&e5&e6) | (e0&e2&e3&e4&e5&~e6) | (~e0&~e1&~e2&~e3&~e4&~e5&e6) | (~e0&~e1&~e2&~e3&e4&~e5&~e6) | (~e0&~e1&~e2&e3&~e4&e5&e6) | (~e0&~e1&~e2&e3&~e4&e5&e6) | (~e0&~e1&~e2&e3&e4&e5&~e6) | (~e0&~e1&~e2&e3&~e4&e5&e6) | (~e0&~e1&e2&~e3&e4&~e5&e6) | (~e0&~e1&e2&e3&~e4&~e5&~e6) | (~e0&~e1&e2&e3&e4&e5&e6) | (~e0&e1&~e2&~e3&~e4&e5&~e6) | (e0&~e1&~e2&~e3&~e4&~e5&~e6));                                                 
	assign b10 = ((e0&e1&~e5&~e6) | (e1&~e2&~e3&e4&~e5&~e6) | (e1&~e2&e3&e4&~e5&e6) | (e1&~e2&e3&e4&e5&~e6) | (e1&e2&~e3&e4&e5&e6) | (e1&e2&e3&~e4&~e5&~e6) | (e0&~e2&e3&~e4&e5&e6) | (e0&~e2&e3&e4&~e5&~e6) | (e0&e2&~e3&e4&~e5&e6) | (e0&e2&~e3&e4&e5&~e6) | (e0&e2&e3&e4&e5&e6) | (~e0&~e1&~e2&~e3&e4&~e5&e6) | (~e0&~e1&~e2&~e3&e4&e5&~e6) | (~e0&~e1&~e2&e3&e4&e5&e6) | (~e0&~e1&e2&~e3&~e4&~e5&~e6) | (~e0&~e1&e2&e3&~e4&~e5&e6) | (~e0&~e1&e2&e3&~e4&e5&~e6) | (~e0&e1&~e2&~e3&~e4&e5&e6) | (e0&~e1&~e2&~e3&~e4&~e5&e6) | (e0&~e1&~e2&~e3&~e4&e5&~e6));                                           
	assign c10 = ((e1&~e2&e3&~e4&e5&~e6) | (e1&e2&~e3&e4&~e5&~e6) | (e1&e2&e3&e4&e5&~e6) | (e0&~e2&e3&~e4&~e5&~e6) | (e0&e2&~e3&~e4&e5&~e6) | (e0&e2&e3&e4&~e5&~e6) | (~e0&~e1&~e2&~e3&~e4&e5&~e6) | (~e0&~e1&~e2&e3&e4&~e5&~e6) | (~e0&~e1&e2&~e3&e4&e5&~e6) | (~e0&e1&~e2&~e3&~e4&~e5&~e6));
	assign d10 = ((e0&e1&~e5&e6) | (e1&e3&~e4&~e5&e6) | (e1&e2&e3&~e5&e6) | (e0&~e3&e4&e5&e6) | (~e0&~e1&~e3&~e4&~e5&e6) | (~e1&~e2&~e3&e4&e5&e6) | (~e0&~e1&e3&~e4&e5&e6) | (~e0&~e1&e2&~e3&~e5&e6) | (~e1&e2&~e3&~e4&~e5&e6) | (~e0&~e1&e2&e3&e5&e6) | (~e1&e2&e3&~e4&e5&e6) | (e0&~e1&~e2&~e3&e5&e6) | (e1&~e2&~e3&e4&~e5&e6) | (e1&~e2&e3&e4&~e5&~e6) | (e1&~e2&e3&e4&e5&e6) | (e1&e2&~e3&~e4&e5&e6) | (e1&e2&~e3&e4&e5&~e6) | (e0&~e2&e3&~e4&e5&~e6) | (e0&~e2&e3&e4&~e5&e6) | (e0&e2&~e3&e4&~e5&~e6) | (e0&e2&e3&e4&e5&~e6) | (~e0&~e1&~e2&~e3&e4&~e5&~e6) | (~e0&~e1&~e2&e3&e4&e5&~e6) | (~e0&~e1&e2&e3&~e4&~e5&~e6) | (~e0&e1&~e2&~e3&~e4&e5&~e6) | (e0&~e1&~e2&~e3&~e4&~e5&~e6));
	assign e10 = ((e6) | (e1&~e2&e3&e4&~e5) | (e1&e2&~e3&e4&e5) | (e0&~e2&e3&~e4&e5) | (e0&e2&~e3&e4&~e5) | (e0&e2&e3&e4&e5) | (~e0&~e1&~e2&~e3&e4&~e5) | (~e0&~e1&~e2&e3&e4&e5) | (~e0&~e1&e2&e3&~e4&~e5) | (~e0&e1&~e2&~e3&~e4&e5) | (e0&~e1&~e2&~e3&~e4&~e5));
	assign f10 = ((~e1&~e2&~e3&e5&e6) | (~e1&~e3&e4&e5&e6) | (e1&~e2&~e3&~e5&e6) | (e1&e3&~e4&~e5&e6) | (e1&~e2&e3&~e4&e5) | (e1&~e2&e3&e5&e6) | (e1&e2&~e3&e4&~e5) | (e1&e2&e4&~e5&e6) | (e1&e2&e3&e4&e5) | (e0&~e2&e3&~e4&~e5) | (e0&~e2&e3&~e5&e6) | (e0&e2&~e3&~e4&e6) | (e0&e2&~e3&~e4&e5) | (e0&e2&~e4&e5&e6) | (e0&e2&e3&e4&~e5) | (~e0&~e1&~e2&~e3&~e4&e6) | (~e0&~e1&~e2&~e3&~e4&e5) | (~e0&~e1&e3&~e4&e5&e6) | (~e0&~e1&~e2&e3&e4&~e5) | (~e0&~e1&e2&~e3&~e5&e6) | (~e0&~e1&e2&~e3&~e5&e6) | (~e0&~e1&e2&~e3&e4&e5) | (~e0&~e1&e2&e4&e5&e6) | (~e0&e1&~e2&~e3&~e4&~e5) | (e1&e2&~e3&~e4&e5&e6));
	assign g10 = ((e0&e1&~e5&e6) | (e1&~e2&e3&~e4&~e5) | (e1&e3&~e4&~e5&e6) | (e1&e2&~e3&~e4&e5) | (e1&e2&e3&e4&~e5) | (e0&~e2&~e3&e4&e5) | (e0&~e3&e4&e5&e6) | (e0&e2&~e3&~e4&~e5) | (e0&e2&e3&~e4&e5) | (~e0&~e1&~e2&~e3&~e4&~e5) | (~e0&~e1&~e3&~e4&~e5&e6) | (~e1&~e2&~e3&e4&e5&e6) | (~e0&~e1&~e2&e3&~e4&e5) | (~e0&~e1&e3&~e4&e5&e6) | (~e0&~e1&e2&~e3&e4&~e5) | (~e0&~e1&e2&e3&e4&e5) | (e0&~e1&~e2&~e3&e5&e6) | (e1&~e2&~e3&e4&~e5&e6) | (e1&~e2&e3&e4&e5&e6) | (e0&~e2&e3&e4&~e5&e6));
endmodule 